-- Team Number 7
-- Vishal Mansuria, Sean McCray 
-- vpm5113@psu.edu, smm7442@psu.edu
-- my_genpulse.vhd
-- Version 1.0 , 10/15/2020
---------------------------------------------------------------------------
-- This VHDL file was developed by Daniel Llamocca (2013).  It may be
-- freely copied and/or distributed at no cost.  Any persons using this
-- file for any purpose do so at their own risk, and are responsible for
-- the results of such use.  Daniel Llamocca does not guarantee that
-- this file is complete, correct, or fit for any particular purpose.
-- NO WARRANTY OF ANY KIND IS EXPRESSED OR IMPLIED.  This notice must
-- accompany any copy of this file.
--------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
--use ieee.math_real.log2;
--use ieee.math_real.ceil;

entity my_genpulse is
	--generic (COUNT: INTEGER:= (10**8)/2); -- (10**8)/2 cycles of T = 10 ns --> 0.5 s
	generic (COUNT: INTEGER:= (10**2)/2 ); -- (10**2)/2 cycles of T = 10 ns --> 0.5us
	port (clock, resetn, E: in std_logic;
			Q: out std_logic_vector ( 31 downto 0);
			z: out std_logic);
end my_genpulse;

architecture Behavioral of my_genpulse is
	constant nbits: INTEGER:= 32;
	signal Qt: std_logic_vector (nbits -1 downto 0);
begin

	process (resetn, clock)
	begin
		if resetn = '0' then
			Qt <= (others => '0');
		elsif (clock'event and clock = '1') then
			if E = '1' then
				if Qt = conv_std_logic_vector (COUNT-1,nbits) then
					Qt <= (others => '0');
				else
					Qt <= Qt + conv_std_logic_vector (1,nbits);
				end if;
			end if;
		end if;
	end process;
	
	z <= '1' when Qt = conv_std_logic_vector (COUNT-1,nbits) else '0';
   Q <= Qt;
	
end Behavioral;

